package types;

/* Example chip-wide parameters */
parameter int NUM_DATA_INPUT_PINS = 8;
parameter int NUM_DATA_OUTPUT_PINS = 4;

/* Put any other shared variables/parameters you want in here. This is automatically available in other modules within the hardware folder! */

endpackage
